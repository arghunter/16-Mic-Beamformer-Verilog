module big_adder(
    input [23:0] in_0,
    input [23:0] in_1,
    input [23:0] in_2,
    input [23:0] in_3,
    input [23:0] in_4,
    input [23:0] in_5,
    input [23:0] in_6,
    input [23:0] in_7,
    input [23:0] in_8,
    output [21:0] sum,
);